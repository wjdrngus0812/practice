module counter (
    input clk,
    input rst_n,
    output reg [3:0] count
);
// TODO: 로직 구현하기
endmodule